library verilog;
use verilog.vl_types.all;
entity testdata is
end testdata;
