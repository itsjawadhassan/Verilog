library verilog;
use verilog.vl_types.all;
entity testmyha is
end testmyha;
