library verilog;
use verilog.vl_types.all;
entity bitwisetest is
end bitwisetest;
