library verilog;
use verilog.vl_types.all;
entity logical_operators is
end logical_operators;
