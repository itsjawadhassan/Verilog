module myand (in1,in2,o);
input in1,in2;
output o;
and a(o,in1,in2);
endmodule

