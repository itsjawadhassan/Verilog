library verilog;
use verilog.vl_types.all;
entity testlogical is
end testlogical;
