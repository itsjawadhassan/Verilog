library verilog;
use verilog.vl_types.all;
entity operatortest is
end operatortest;
