library verilog;
use verilog.vl_types.all;
entity testcircuit is
end testcircuit;
