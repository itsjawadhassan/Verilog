library verilog;
use verilog.vl_types.all;
entity testgate is
end testgate;
